-- Dimitris Tsiompikas 3180223
-- Antwnhs Detshs 3190054
-- Petros Tsotsi 3180193


LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY MUX8_1_16BIT IS

PORT (IN0,IN1,IN2,IN3,IN4,IN5,IN6,IN7 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		SEL : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		OUT1 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
		
		
END MUX8_1_16BIT;


ARCHITECTURE logic_structural OF MUX8_1_16BIT IS

COMPONENT MUX8_1 IS

PORT (IN0,IN1,IN2,IN3,IN4,IN5,IN6,IN7 : IN STD_LOGIC;
		SEL : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		OUT1 : OUT STD_LOGIC);
		
		
END COMPONENT;

BEGIN

	V0 : MUX8_1 port map (IN0(0),IN1(0),IN2(0),IN3(0),IN4(0),IN5(0),IN6(0),IN7(0),SEL,OUT1(0)); 
	V1 : MUX8_1 port map (IN0(1),IN1(1),IN2(1),IN3(1),IN4(1),IN5(1),IN6(1),IN7(1),SEL,OUT1(1));
	V2 : MUX8_1 port map (IN0(2),IN1(2),IN2(2),IN3(2),IN4(2),IN5(2),IN6(2),IN7(2),SEL,OUT1(2));
	V3 : MUX8_1 port map (IN0(3),IN1(3),IN2(3),IN3(3),IN4(3),IN5(3),IN6(3),IN7(3),SEL,OUT1(3));
	V4 : MUX8_1 port map (IN0(4),IN1(4),IN2(4),IN3(4),IN4(4),IN5(4),IN6(4),IN7(4),SEL,OUT1(4));
	V5 : MUX8_1 port map (IN0(5),IN1(5),IN2(5),IN3(5),IN4(5),IN5(5),IN6(5),IN7(5),SEL,OUT1(5));
	V6 : MUX8_1 port map (IN0(6),IN1(6),IN2(6),IN3(6),IN4(6),IN5(6),IN6(6),IN7(6),SEL,OUT1(6));
	V7 : MUX8_1 port map (IN0(7),IN1(7),IN2(7),IN3(7),IN4(7),IN5(7),IN6(7),IN7(7),SEL,OUT1(7));
	V8 : MUX8_1 port map (IN0(8),IN1(8),IN2(8),IN3(8),IN4(8),IN5(8),IN6(8),IN7(8),SEL,OUT1(8));
	V9 : MUX8_1 port map (IN0(9),IN1(9),IN2(9),IN3(9),IN4(9),IN5(9),IN6(9),IN7(9),SEL,OUT1(9));
	V10 : MUX8_1 port map (IN0(10),IN1(10),IN2(10),IN3(10),IN4(10),IN5(10),IN6(10),IN7(10),SEL,OUT1(10));
	V11 : MUX8_1 port map (IN0(11),IN1(11),IN2(11),IN3(11),IN4(11),IN5(11),IN6(11),IN7(11),SEL,OUT1(11));
	V12 : MUX8_1 port map (IN0(12),IN1(12),IN2(12),IN3(12),IN4(12),IN5(12),IN6(12),IN7(12),SEL,OUT1(12));
	V13 : MUX8_1 port map (IN0(13),IN1(13),IN2(13),IN3(13),IN4(13),IN5(13),IN6(13),IN7(13),SEL,OUT1(13));
	V14 : MUX8_1 port map (IN0(14),IN1(14),IN2(14),IN3(14),IN4(14),IN5(14),IN6(14),IN7(14),SEL,OUT1(14));
	V15 : MUX8_1 port map (IN0(15),IN1(15),IN2(15),IN3(15),IN4(15),IN5(15),IN6(15),IN7(15),SEL,OUT1(15));
	
END logic_structural;