-- Dimitris Tsiompikas 3180223
-- Antwnhs Detshs 3190054
-- Petros Tsotsi 3180193


LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY OR_3 IS 

PORT ( IN1, IN2, IN3 : IN STD_LOGIC;
		 OUT1 : OUT STD_LOGIC);
		 
END OR_3;


ARCHITECTURE LOGICFUNC OF OR_3 IS

COMPONENT OR_2 IS
PORT ( IN1, IN2 : IN STD_LOGIC;
		 OUT1 : OUT STD_LOGIC);
		
END COMPONENT;
	signal C : std_logic;
BEGIN 
	V0 : OR_2 port map (IN1,IN2,C);
	V1 : OR_2 port map (C,IN3,OUT1);
	
END LOGICFUNC;