-- Dimitris Tsiompikas 3180223
-- Antwnhs Detshs 3190054
-- Petros Tsotsi 3180193


LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;



ENTITY MUX8_1 IS

PORT (IN0,IN1,IN2,IN3,IN4,IN5,IN6,IN7 : IN STD_LOGIC;
		SEL : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		OUT1 : OUT STD_LOGIC);
		
		
END MUX8_1;


ARCHITECTURE LOGICFUNC OF MUX8_1 IS


COMPONENT NOT1 IS 

PORT ( A : IN STD_LOGIC;
		 Q : OUT STD_LOGIC);
		 
END COMPONENT;



COMPONENT AND_4 IS 

PORT ( IN1 , IN2, IN3, IN4 : IN STD_LOGIC;
		 OUT1 : OUT STD_LOGIC);
		 
END COMPONENT;



COMPONENT OR_8 IS 

PORT ( IN1, IN2, IN3, IN4 , IN5 , IN6 , IN7, IN8 : IN STD_LOGIC;
		 OUT1 : OUT STD_LOGIC);
		 
END COMPONENT;



SIGNAL NOTSEL : STD_LOGIC_VECTOR(2 DOWNTO 0);

SIGNAL S0,S1,S2,S3,S4,S5,S6,S7 : STD_LOGIC;


BEGIN

-- NOT GATE FOR SELECTOR BITS

V0: NOT1 PORT MAP (SEL(0) , NOTSEL(0));
V1: NOT1 PORT MAP (SEL(1) , NOTSEL(1));
V2: NOT1 PORT MAP (SEL(2) , NOTSEL(2));



-- IF OPCODE IS '000' , SELECT IN1 

V3: AND_4 PORT MAP (NOTSEL(2) , NOTSEL(1) , NOTSEL(0) , IN0 , S0);


-- IF OPCODE IS '001' , SELECT IN2 

V4: AND_4 PORT MAP (NOTSEL(2) , NOTSEL(1) , SEL(0) , IN1, S1);


-- IF OPCODE IS '010' , SELECT IN3

V5: AND_4 PORT MAP (NOTSEL(2), SEL(1) , NOTSEL(0) , IN2, S2);


-- IF OPCODE IS '011' , SELECT IN4 

V6: AND_4 PORT MAP (NOTSEL(2) , SEL(1) , SEL(0) , IN3 , S3);


-- IF OPCODE IS '100' , SELECT IN5

V7: AND_4 PORT MAP (SEL(2) , NOTSEL(1) , NOTSEL(0), IN4, S4);


-- IF OPCODE IS '101' , SELECT IN6 

V8: AND_4 PORT MAP (SEL(2) , NOTSEL(1) , SEL(0) , IN5 , S5);


-- IF OPCODE IS '110' , SELECT IN7 

V9: AND_4 PORT MAP (SEL(2) , SEL(1) , NOTSEL(0) , IN6 , S6);


-- IF OPCODE IS '111' , SELECT IN8 


V10: AND_4 PORT MAP (SEL(2) , SEL(1), SEL(0) , IN7 , S7);


-- FINAL MULTIPLEXER OUTPUT

V11: OR_8 PORT MAP (S0,S1,S2,S3,S4,S5,S6,S7 , OUT1 );




END LOGICFUNC;