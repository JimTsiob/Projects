-- Dimitris Tsiompikas 3180223
-- Antwnhs Detshs 3190054
-- Petros Tsotsi 3180193


LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY AND_2 IS 

PORT ( IN1 , IN2 : IN STD_LOGIC;
		 OUT1 : OUT STD_LOGIC);
		 
END AND_2;



ARCHITECTURE LOGICFUNC OF AND_2 IS

BEGIN 

	OUT1 <= IN1 AND IN2;
	
END LOGICFUNC;

