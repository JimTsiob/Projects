-- Dimitrios Tsiompikas 3180223
-- Antonis Detsis 3190054
-- Petros Tsotsi 3180193

LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY DEC_3_TO_8 IS
PORT(
		Input : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		Output : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
);
END DEC_3_TO_8;

ARCHITECTURE LogicFunc OF DEC_3_TO_8 IS
BEGIN
	WITH Input SELECT
		Output <= "00000001" WHEN "000",
					 "00000010" WHEN "001",
					 "00000100" WHEN "010",
					 "00001000" WHEN "011",
					 "00010000" WHEN "100",
					 "00100000" WHEN "101",
					 "01000000" WHEN "110",
					 "10000000" WHEN "111",
					 "00000000" WHEN OTHERS;

END LogicFunc;