-- Dimitris Tsiompikas 3180223
-- Antwnhs Detshs 3190054
-- Petros Tsotsi 3180193


LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY XOR_3 IS 

PORT ( IN1, IN2, IN3 : IN STD_LOGIC;
		 OUT1 : OUT STD_LOGIC);
		 
END XOR_3;


ARCHITECTURE LOGICFUNC OF XOR_3 IS

COMPONENT XOR_2 IS

PORT ( A ,B : IN STD_LOGIC ;
		 Z : OUT STD_LOGIC);
		 
END COMPONENT;

signal C : std_logic;

BEGIN 
	V0 : XOR_2 PORT MAP (IN1,IN2,C);
	V1 : XOR_2 PORT MAP (C,IN3,OUT1);
	
	
END LOGICFUNC;